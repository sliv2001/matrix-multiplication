
module unsaved (
	clk_clk,
	reset_reset_n,
	onchip_memory2_0_reset1_reset,
	onchip_memory2_0_reset1_reset_req);	

	input		clk_clk;
	input		reset_reset_n;
	input		onchip_memory2_0_reset1_reset;
	input		onchip_memory2_0_reset1_reset_req;
endmodule
